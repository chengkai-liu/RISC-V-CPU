`include "defines.v"

module mctrl(
    input wire              rst,
    input wire              rdy,
    
);

endmodule // mctrl