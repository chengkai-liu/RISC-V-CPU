`include "defines.v"
//todo no need
module mctrl(
    input wire                  rst,
    input wire                  rdy,
    
    // from if
    input wire                  if_mctrl_req_i,
    // from mem for load/store
    input wire                  mem_mctrl_req_i,

    input wire                  
);

endmodule // mctrl