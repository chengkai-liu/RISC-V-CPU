`include "defines.v"

module icache(
    input wire              clk,
    input wire              rst,
    input wire              rdy,

);

endmodule // icache