`include "defines.v"

module ctrl(
    
);

endmodule // ctrl