`include "defines.v"

module dcache(
    
);

endmodule // dcache