`include "defines.v"

module if(
    input wire rst,


);

endmodule // if